* G:\ESIMworkplace\hack\hack.cir

* EESchema Netlist Version 1.1 (Spice format) creation date: 11/07/24 00:59:16

* To exclude a component from the Spice Netlist add [Spice_Netlist_Enabled] user FIELD set to: N
* To reorder the component spice node sequence add [Spice_Node_Sequence] user FIELD and define sequence: 2,1,0

* Sheet Name: /
scmode1  SKY130mode		
SC2  Net-_SC1-Pad1_ A GND GND sky130_fd_pr__nfet_01v8		
SC1  Net-_SC1-Pad1_ A Net-_SC1-Pad3_ Net-_SC1-Pad3_ sky130_fd_pr__pfet_01v8		
SC3  CARRY A Net-_SC1-Pad3_ Net-_SC1-Pad3_ sky130_fd_pr__pfet_01v8		
SC5  SUM C A Net-_SC1-Pad3_ sky130_fd_pr__pfet_01v8		
SC4  CARRY A C GND sky130_fd_pr__nfet_01v8		
SC6  SUM C Net-_SC1-Pad1_ GND sky130_fd_pr__nfet_01v8		
v1  A GND pulse		
v2  C GND pulse		
U1  A plot_v1		
U2  C plot_v1		
U4  SUM plot_v1		
U3  CARRY plot_v1		
v3  Net-_SC1-Pad3_ GND DC		
SC7  SUM GND sky130_fd_pr__cap_mim_m3_1		

.end
